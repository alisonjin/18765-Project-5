`timescale 1ns / 1ps

module nm_testbench();

   reg CK, scan_en, bist_en, TPG_reset, COMP_reset, SI_chain1, SI_chain2, SI_chain3, SI_chain4, SI_chain5, SI_chain6, SI_chain7, 
   SO_chain1, SO_chain2, SO_chain3, SO_chain4, SO_chain5, SO_chain6, SO_chain7;  // Add new pins in your design
   reg [246:0] LFSR;
   wire [249:0] TEST_OUT;
   wire g89,g94,g98,g102,g107,g301,g306,g310,g314,g319,g557,g558,g559,g560,g561,g562,g563,g564,g705,g639,g567,g45,g42,g39,g702,g32,g38,g46,g36,g47,g40,g37,g41,g22,g44,g23;
   wire g2584_orig,g3222_orig,g3600_orig,g4307_orig,g4321_orig,g4422_orig,g4809_orig,g5137_orig,g5468_orig,g5469_orig,g5692_orig,g6282_orig,g6284_orig,g6360_orig,g6362_orig,g6364_orig,g6366_orig,g6368_orig,g6370_orig,g6372_orig,g6374_orig,g6728_orig,g1290_orig,g4121_orig,g4108_orig,g4106_orig,g4103_orig,g1293_orig,g4099_orig,g4102_orig,g4109_orig,g4100_orig,g4112_orig,g4105_orig,g4101_orig,g4110_orig,g4104_orig,g4107_orig,g4098_orig;
   wire g2584,g3222,g3600,g4307,g4321,g4422,g4809,g5137,g5468,g5469,g5692,g6282,g6284,g6360,g6362,g6364,g6366,g6368,g6370,g6372,g6374,g6728,g1290,g4121,g4108,g4106,g4103,g1293,g4099,g4102,g4109,g4100,g4112,g4105,g4101,g4110,g4104,g4107,g4098;
   integer f, i;

    // combination circuit
    s9234_comb comb(g89,g94,g98,g102,g107,g301,g306,g310,g314,g319,g557,g558,g559,g560,g561,
        g562,g563,g564,g705,g639,g567,g45,g42,g39,g702,g32,g38,g46,g36,g47,g40,g37,
        g41,g22,g44,g23, 
        
        g678,g332,g123,g207,g695,g461,g18, g292,g331,g689,g24, g465,g84, g291,g676,g622,g117,g278,g128,g598,g554,g496,g179,g48, g590,g551,g682,g11, g606,g188,g646,g327,g361,g289,g398,g684,g619,g208,g248,g390,g625,g681,g437,g276,g3,  g323,g224,g685,g43, g157,g282,g697,g206,g449,g118,g528,g284,g426,g634,g669,g520,g281,g175,g15, g631,g69, g693,g337,g457,g486,g471,g328,g285,g418,g402,g297,g212,g410,g430,g33, g662,g453,g269,g574,g441,g664,g349,g211,g586,g571,g29, g326,g698,g654,g293,g690,g445,g374,g6,  g687,g357,g386,g504,g665,g166,g541,g74, g338,g696,g516,g536,g683,g353,g545,g254,g341,g290,g2,  g287,g336,g345,g628,g679,g28, g688,g283,g613,g10, g14, g680,g143,g672,g667,g366,g279,g492,g170,g686,g288,g638,g602,g642,g280,g663,g610,g148,g209,g675,g478,g122,g54, g594,g286,g489,g616,g79, g218,g242,g578,g184,g119,g668,g139,g422,g210,g394,g230,g25, g204,g658,g650,g378,g508,g548,g370,g406,g236,g500,g205,g197,g666,g114,g524,g260,g111,g131,g7,  g19, g677,g582,g485,g699,g193,g135,g382,g414,g434,g266,g49, g152,g692,g277,g127,g161,g512,g532,g64, g694,g691,g1,g59,
        
        g2584,g3222,g3600,g4307,g4321,g4422,g4809,g5137,g5468,g5469,g5692,g6282,
        g6284,g6360,g6362,g6364,g6366,g6368,g6370,g6372,g6374,g6728,g1290,g4121,
        g4108,g4106,g4103,g1293,g4099,g4102,g4109,g4100,g4112,g4105,g4101,g4110,
        g4104,g4107,g4098,
        
        g4130,g6823,g6940,g6102,g4147,g4841,g6725,g3232,g4119,g4141,g6726,g6507,g6590,g3231,g5330,g5147,g4839,g6105,g5138,g4122,g6827,g6745,g6405,g6729,g6595,g6826,g4134,g6599,g4857,g6406,g5148,g4117,g6582,g3229,g5700,g4136,g4858,g5876,g3239,g5698,g5328,g4133,g4847,g5877,g6597,g4120,g3235,g4137,g6407,g5470,g6841,g4149,g6101,g4844,g4113,g6504,g3224,g4855,g4424,g5582,g6502,g6107,g5472,g6602,g5581,g6587,g4145,g2585,g4842,g2586,g1291,g4118,g3225,g4853,g4849,g6512,g3233,g4851,g4856,g6854,g1831,g4843,g6510,g6591,g4846,g1288,g5478,g6840,g6594,g5580,g6853,g4840,g4150,g5490,g6511,g4142,g4845,g5694,g6722,g4139,g5480,g5697,g6498,g4126,g5471,g6505,g6588,g5475,g4148,g6501,g6506,g4135,g5479,g6824,g3240,g5476,g3230,g6721,g3227,g6925,g5477,g5489,g4131,g6727,g4140,g6842,g4423,g6723,g6724,g4132,g6401,g5491,g4127,g6278,g6106,g6744,g6404,g4138,g3228,g1289,g4123,g4658,g5878,g4125,g4124,g5874,g6103,g1294,g1292,g4115,g6584,g6596,g3226,g2587,g4657,g6589,g3234,g3238,g6592,g5473,g4114,g6800,g5141,g4854,g6839,g5699,g3236,g6601,g5875,g4425,g5329,g5695,g6499,g6825,g5693,g4850,g3237,g6497,g6100,g6509,g4128,g4116,g6503,g3241,g6277,g5139,g6598,g6600,g4129,g6593,g6801,g4426,g5474,g5140,g5696,g4852,g4848,g4659,g6583,g6402,g4144,g6104,g6941,g6403,g6500,g6508,g6586,g4146,g4143,g6720,g6585
    );
   
   // regular PI
   assign {g89,g94,g98,g102,g107,g301,g306,g310,g314,g319,g557,g558,g559,g560,g561,g562,g563,g564,g705,g639,g567,g45,g42,g39,g702,g32,g38,g46,g36,g47,g40,g37,g41,g22,g44,g23} = LFSR[246:211];
   
   // DFF inputs
   assign {g678,g332,g123,g207,g695,g461,g18, g292,g331,g689,g24, g465,g84, g291,
   g676,g622,g117,g278,g128,g598,g554,g496,g179,g48, g590,g551,g682,g11, g606,g188,
   g646,g327,g361,g289,g398,g684,g619,g208,g248,g390,g625,g681,g437,g276,g3,  g323,
   g224,g685,g43, g157,g282,g697,g206,g449,g118,g528,g284,g426,g634,g669,g520,g281,
   g175,g15, g631,g69, g693,g337,g457,g486,g471,g328,g285,g418,g402,g297,g212,g410,
   g430,g33, g662,g453,g269,g574,g441,g664,g349,g211,g586,g571,g29, g326,g698,g654,
   g293,g690,g445,g374,g6,  g687,g357,g386,g504,g665,g166,g541,g74, g338,g696,g516,
   g536,g683,g353,g545,g254,g341,g290,g2,  g287,g336,g345,g628,g679,g28, g688,g283,
   g613,g10, g14, g680,g143,g672,g667,g366,g279,g492,g170,g686,g288,g638,g602,g642,
   g280,g663,g610,g148,g209,g675,g478,g122,g54, g594,g286,g489,g616,g79, g218,g242,
   g578,g184,g119,g668,g139,g422,g210,g394,g230,g25, g204,g658,g650,g378,g508,g548,
   g370,g406,g236,g500,g205,g197,g666,g114,g524,g260,g111,g131,g7,  g19, g677,g582,
   g485,g699,g193,g135,g382,g414,g434,g266,g49, g152,g692,g277,g127,g161,g512,g532,
   g64, g694,g691,g1,  g59} = LFSR[210:0];

   assign TEST_OUT[249:0] = {g2584,g3222,g3600,g4307,g4321,g4422,g4809,g5137,g5468,
   g5469,g5692,g6282,g6284,g6360,g6362,g6364,g6366,g6368,g6370,g6372,g6374,g6728,g1290,
   g4121,g4108,g4106,g4103,g1293,g4099,g4102,g4109,g4100,g4112,g4105,g4101,g4110,g4104,
   g4107,g4098,g4130,g6823,g6940,g6102,g4147,g4841,g6725,g3232,g4119,g4141,g6726,g6507,
   g6590,g3231,g5330,g5147,g4839,g6105,g5138,g4122,g6827,g6745,g6405,g6729,g6595,g6826,
   g4134,g6599,g4857,g6406,g5148,g4117,g6582,g3229,g5700,g4136,g4858,g5876,g3239,g5698,
   g5328,g4133,g4847,g5877,g6597,g4120,g3235,g4137,g6407,g5470,g6841,g4149,g6101,g4844,
   g4113,g6504,g3224,g4855,g4424,g5582,g6502,g6107,g5472,g6602,g5581,g6587,g4145,g2585,
   g4842,g2586,g1291,g4118,g3225,g4853,g4849,g6512,g3233,g4851,g4856,g6854,g1831,g4843,
   g6510,g6591,g4846,g1288,g5478,g6840,g6594,g5580,g6853,g4840,g4150,g5490,g6511,g4142,
   g4845,g5694,g6722,g4139,g5480,g5697,g6498,g4126,g5471,g6505,g6588,g5475,g4148,g6501,
   g6506,g4135,g5479,g6824,g3240,g5476,g3230,g6721,g3227,g6925,g5477,g5489,g4131,g6727,
   g4140,g6842,g4423,g6723,g6724,g4132,g6401,g5491,g4127,g6278,g6106,g6744,g6404,g4138,
   g3228,g1289,g4123,g4658,g5878,g4125,g4124,g5874,g6103,g1294,g1292,g4115,g6584,g6596,
   g3226,g2587,g4657,g6589,g3234,g3238,g6592,g5473,g4114,g6800,g5141,g4854,g6839,g5699,
   g3236,g6601,g5875,g4425,g5329,g5695,g6499,g6825,g5693,g4850,g3237,g6497,g6100,g6509,
   g4128,g4116,g6503,g3241,g6277,g5139,g6598,g6600,g4129,g6593,g6801,g4426,g5474,g5140,
   g5696,g4852,g4848,g4659,g6583,g6402,g4144,g6104,g6941,g6403,g6500,g6508,g6586,g4146,
   g4143,g6720,g6585};


   initial begin
      f = $fopen("output.txt","w");
      CK=0;
      scan_en=0;  // Configure the pins in your design
      bist_en=1;
      TPG_reset=1;
      COMP_reset=0;
    //   scan_in=0;

      SI_chain1 = 0;
      SI_chain2 = 0;
      SI_chain3 = 0;
      SI_chain4 = 0;
      SI_chain5 = 0;
      SI_chain6 = 0;
      SI_chain7 = 0;
      #20;

#5 CK=0;
#5 LFSR=247'b100000011111110101010011001110111010000001000000111111101010100110011101110100000010000001111111010101001100111011100000000100000011111110101010011001110111000000001000000111111101010100110011101100000000010000001111111010101001100111010000000000011111110101010011001110111010000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b010110001101111011010110110010010001000000101100011011110110101101100100100000000001011000110111101101011011001001000000010010110001101111011010110110010010000000100101100011011110110101101100100100000101001011000110111101101011011001000000010110001101111011010110110010010001100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b110000101111100101011100110100010011000001100001011111001010111001101000100100000111000010111110010101110011010001000000001110000101111100101011100110100010000000011100001011111001010111001101000100000000111000010111110010101110011010000000010000101111100101011100110100010011100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b110001010000110000010000001111111010000001100010100001100000100000011111110100000111000101000011000001000000111111100000011110001010000110000010000001111111000000111100010100001100000100000011111100000001111000101000011000001000000111110000010001010000110000010000001111111010100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b101001100111011101001011000110111101000001010011001110111010010110001101111000000010100110011101110100101100011011110000010101001100111011101001011000110111000000101010011001110111010010110001101100000101010100110011101110100101100011010000001001100111011101001011000110111101100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b101011011001001000111000010111110010000001010110110010010001110000101111100100000110101101100100100011100001011111000000001101011011001001000111000010111110000001011010110110010010001110000101111100000110110101101100100100011100001011110000001011011001001000111000010111110010100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b101110011010001001111000101000011000000001011100110100010011110001010000110000000010111001101000100111100010100001100000010101110011010001001111000101000011000000101011100110100010011110001010000100000001010111001101000100111100010100000000001110011010001001111000101000011000000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b001000000111111101010100110011101110000000010000001111111010101001100111011100000000100000011111110101010011001110110000000001000000111111101010100110011101000000000010000001111111010101001100111000000100000100000011111110101010011001110000001000000111111101010100110011101110100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b100101100011011110110101101100100100000001001011000110111101101011011001001000000010010110001101111011010110110010010000010100101100011011110110101101100100000001101001011000110111101101011011001000000111010010110001101111011010110110010000000101100011011110110101101100100100000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b011100001011111001010111001101000100000000111000010111110010101110011010001000000001110000101111100101011100110100010000000011100001011111001010111001101000000001000111000010111110010101110011010000000010001110000101111100101011100110100000011100001011111001010111001101000100100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b111100010100001100000100000011111110000001111000101000011000001000000111111100000011110001010000110000010000001111110000000111100010100001100000100000011111000001001111000101000011000001000000111100000010011110001010000110000010000001110000011100010100001100000100000011111110100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b101010011001110111010010110001101111000001010100110011101110100101100011011100000010101001100111011101001011000110110000010101010011001110111010010110001101000001101010100110011101110100101100011000000111010101001100111011101001011000110000001010011001110111010010110001101111000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b011010110110010010001110000101111100000000110101101100100100011100001011111000000101101011011001001000111000010111110000011011010110110010010001110000101111000001110110101101100100100011100001011100000111101101011011001001000111000010110000011010110110010010001110000101111100100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b101011100110100010011110001010000110000001010111001101000100111100010100001100000010101110011010001001111000101000010000000101011100110100010011110001010000000001001010111001101000100111100010100000000110010101110011010001001111000101000000001011100110100010011110001010000110000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b000010000001111111010101001100111011000000000100000011111110101010011001110100000000001000000111111101010100110011100000010000010000001111111010101001100111000001100000100000011111110101010011001100000011000001000000111111101010100110010000000010000001111111010101001100111011100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b101001011000110111101101011011001001000001010010110001101111011010110110010000000110100101100011011110110101101100100000011101001011000110111101101011011001000000111010010110001101111011010110110000000101110100101100011011110110101101100000001001011000110111101101011011001001000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b000111000010111110010101110011010001000000001110000101111100101011100110100000000100011100001011111001010111001101000000001000111000010111110010101110011010000000010001110000101111100101011100110100000100100011100001011111001010111001100000000111000010111110010101110011010001000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b001111000101000011000001000000111111000000011110001010000110000010000001111100000100111100010100001100000100000011110000001001111000101000011000001000000111000000010011110001010000110000010000001100000000100111100010100001100000100000010000001111000101000011000001000000111111100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b101010100110011101110100101100011011000001010101001100111011101001011000110100000110101010011001110111010010110001100000011101010100110011101110100101100011000001111010101001100111011101001011000100000111110101010011001110111010010110000000001010100110011101110100101100011011100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b110110101101100100100011100001011111000001101101011011001001000111000010111100000111011010110110010010001110000101110000011110110101101100100100011100001011000000111101101011011001001000111000010100000101111011010110110010010001110000100000010110101101100100100011100001011111000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b001010111001101000100111100010100001000000010101110011010001001111000101000000000100101011100110100010011110001010000000011001010111001101000100111100010100000001110010101110011010001001111000101000000111100101011100110100010011110001010000001010111001101000100111100010100001100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b100000100000011111110101010011001110000001000001000000111111101010100110011100000110000010000001111111010101001100110000001100000100000011111110101010011001000000011000001000000111111101010100110000000000110000010000001111111010101001100000000000100000011111110101010011001110100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b111010010110001101111011010110110010000001110100101100011011110110101101100100000011101001011000110111101101011011000000010111010010110001101111011010110110000001101110100101100011011110110101101100000111011101001011000110111101101011010000011010010110001101111011010110110010000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b010001110000101111100101011100110100000000100011100001011111001010111001101000000001000111000010111110010101110011010000010010001110000101111100101011100110000000100100011100001011111001010111001100000001001000111000010111110010101110010000010001110000101111100101011100110100000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b010011110001010000110000010000001111000000100111100010100001100000100000011100000001001111000101000011000001000000110000000010011110001010000110000010000001000001000100111100010100001100000100000000000010001001111000101000011000001000000000010011110001010000110000010000001111100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b111010101001100111011101001011000110000001110101010011001110111010010110001100000111101010100110011101110100101100010000011111010101001100111011101001011000000001111110101010011001110111010010110000000111111101010100110011101110100101100000011010101001100111011101001011000110100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b111101101011011001001000111000010111000001111011010110110010010001110000101100000011110110101101100100100011100001010000010111101101011011001001000111000010000001101111011010110110010010001110000100000011011110110101101100100100011100000000011101101011011001001000111000010111100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b110010101110011010001001111000101000000001100101011100110100010011110001010000000111001010111001101000100111100010100000011110010101110011010001001111000101000001111100101011100110100010011110001000000011111001010111001101000100111100010000010010101110011010001001111000101000000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b011000001000000111111101010100110011000000110000010000001111111010101001100100000001100000100000011111110101010011000000000011000001000000111111101010100110000000000110000010000001111111010101001100000100001100000100000011111110101010010000011000001000000111111101010100110011100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b101110100101100011011110110101101100000001011101001011000110111101101011011000000110111010010110001101111011010110110000011101110100101100011011110110101101000000111011101001011000110111101101011000000001110111010010110001101111011010110000001110100101100011011110110101101100100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b100100011100001011111001010111001101000001001000111000010111110010101110011000000010010001110000101111100101011100110000000100100011100001011111001010111001000001001001000111000010111110010101110000000110010010001110000101111100101011100000000100011100001011111001010111001101000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b000100111100010100001100000100000011000000001001111000101000011000001000000100000100010011110001010000110000010000000000001000100111100010100001100000100000000001010001001111000101000011000001000000000110100010011110001010000110000010000000000100111100010100001100000100000011100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b111110101010011001110111010010110001000001111101010100110011101110100101100000000111111010101001100111011101001011000000011111110101010011001110111010010110000000111111101010100110011101110100101100000001111111010101001100111011101001010000011110101010011001110111010010110001100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b101111011010110110010010001110000101000001011110110101101100100100011100001000000110111101101011011001001000111000010000001101111011010110110010010001110000000000011011110110101101100100100011100000000000110111101101011011001001000111000000001111011010110110010010001110000101100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b111100101011100110100010011110001010000001111001010111001101000100111100010100000111110010101110011010001001111000100000001111100101011100110100010011110001000001011111001010111001101000100111100000000010111110010101110011010001001111000000011100101011100110100010011110001010000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b000110000010000001111111010101001100000000001100000100000011111110101010011000000000011000001000000111111101010100110000010000110000010000001111111010101001000000100001100000100000011111110101010000000101000011000001000000111111101010100000000110000010000001111111010101001100100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b111011101001011000110111101101011011000001110111010010110001101111011010110100000011101110100101100011011110110101100000000111011101001011000110111101101011000001001110111010010110001101111011010100000110011101110100101100011011110110100000011011101001011000110111101101011011000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b001001000111000010111110010101110011000000010010001110000101111100101011100100000100100100011100001011111001010111000000011001001000111000010111110010101110000000110010010001110000101111100101011100000101100100100011100001011111001010110000001001000111000010111110010101110011000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b010001001111000101000011000001000000000000100010011110001010000110000010000000000101000100111100010100001100000100000000011010001001111000101000011000001000000000110100010011110001010000110000010000000001101000100111100010100001100000100000010001001111000101000011000001000000100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b111111101010100110011101110100101100000001111111010101001100111011101001011000000011111110101010011001110111010010110000000111111101010100110011101110100101000000001111111010101001100111011101001000000000011111110101010011001110111010010000011111101010100110011101110100101100000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b011011110110101101100100100011100001000000110111101101011011001001000111000000000001101111011010110110010010001110000000000011011110110101101100100100011100000001000110111101101011011001001000111000000110001101111011010110110010010001110000011011110110101101100100100011100001000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b011111001010111001101000100111100010000000111110010101110011010001001111000100000101111100101011100110100010011110000000001011111001010111001101000100111100000000010111110010101110011010001001111000000000101111100101011100110100010011110000011111001010111001101000100111100010100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b100001100000100000011111110101010011000001000011000001000000111111101010100100000010000110000010000001111111010101000000010100001100000100000011111110101010000000101000011000001000000111111101010100000001010000110000010000001111111010100000000001100000100000011111110101010011000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b001110111010010110001101111011010110000000011101110100101100011011110110101100000100111011101001011000110111101101010000011001110111010010110001101111011010000000110011101110100101100011011110110100000001100111011101001011000110111101100000001110111010010110001101111011010110100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b110010010001110000101111100101011100000001100100100011100001011111001010111000000011001001000111000010111110010101110000010110010010001110000101111100101011000001101100100100011100001011111001010100000011011001001000111000010111110010100000010010010001110000101111100101011100100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b110100010011110001010000110000010000000001101000100111100010100001100000100000000011010001001111000101000011000001000000000110100010011110001010000110000010000001001101000100111100010100001100000100000110011010001001111000101000011000000000010100010011110001010000110000010000000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b001111111010101001100111011101001011000000011111110101010011001110111010010100000000111111101010100110011101110100100000000001111111010101001100111011101001000000000011111110101010011001110111010000000000000111111101010100110011101110100000001111111010101001100111011101001011000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b000110111101101011011001001000111000000000001101111011010110110010010001110000000100011011110110101101100100100011100000011000110111101101011011001001000111000000110001101111011010110110010010001100000101100011011110110101101100100100010000000110111101101011011001001000111000000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b010111110010101110011010001001111000000000101111100101011100110100010011110000000001011111001010111001101000100111100000000010111110010101110011010001001111000000000101111100101011100110100010011100000100001011111001010111001101000100110000010111110010101110011010001001111000100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b101000011000001000000111111101010100000001010000110000010000001111111010101000000010100001100000100000011111110101010000000101000011000001000000111111101010000000001010000110000010000001111111010100000100010100001100000100000011111110100000001000011000001000000111111101010100100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b110011101110100101100011011110110101000001100111011101001011000110111101101000000011001110111010010110001101111011010000000110011101110100101100011011110110000001001100111011101001011000110111101100000010011001110111010010110001101111010000010011101110100101100011011110110101100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b101100100100011100001011111001010111000001011001001000111000010111110010101100000110110010010001110000101111100101010000001101100100100011100001011111001010000001011011001001000111000010111110010100000010110110010010001110000101111100100000001100100100011100001011111001010111000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b001101000100111100010100001100000100000000011010001001111000101000011000001000000100110100010011110001010000110000010000011001101000100111100010100001100000000001110011010001001111000101000011000000000011100110100010011110001010000110000000001101000100111100010100001100000100000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b000011111110101010011001110111010010000000000111111101010100110011101110100100000000001111111010101001100111011101000000000000011111110101010011001110111010000001000000111111101010100110011101110100000010000001111111010101001100111011100000000011111110101010011001110111010010100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b110001101111011010110110010010001110000001100011011110110101101100100100011100000011000110111101101011011001001000110000010110001101111011010110110010010001000000101100011011110110101101100100100000000001011000110111101101011011001001000000010001101111011010110110010010001110000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b000101111100101011100110100010011110000000001011111001010111001101000100111100000000010111110010101110011010001001110000010000101111100101011100110100010011000001100001011111001010111001101000100100000111000010111110010101110011010001000000000101111100101011100110100010011110000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b001010000110000010000001111111010101000000010100001100000100000011111110101000000000101000011000001000000111111101010000010001010000110000010000001111111010000001100010100001100000100000011111110100000111000101000011000001000000111111100000001010000110000010000001111111010101000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b001100111011101001011000110111101101000000011001110111010010110001101111011000000100110011101110100101100011011110110000001001100111011101001011000110111101000001010011001110111010010110001101111000000010100110011101110100101100011011110000001100111011101001011000110111101101000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b011011001001000111000010111110010101000000110110010010001110000101111100101000000101101100100100011100001011111001010000001011011001001000111000010111110010000001010110110010010001110000101111100100000110101101100100100011100001011111000000011011001001000111000010111110010101100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b110011010001001111000101000011000001000001100110100010011110001010000110000000000111001101000100111100010100001100000000001110011010001001111000101000011000000001011100110100010011110001010000110000000010111001101000100111100010100001100000010011010001001111000101000011000001000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b000000111111101010100110011101110100000000000001111111010101001100111011101000000100000011111110101010011001110111010000001000000111111101010100110011101110000000010000001111111010101001100111011100000000100000011111110101010011001110110000000000111111101010100110011101110100100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b101100011011110110101101100100100011000001011000110111101101011011001001000100000010110001101111011010110110010010000000000101100011011110110101101100100100000001001011000110111101101011011001001000000010010110001101111011010110110010010000001100011011110110101101100100100011100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b100001011111001010111001101000100111000001000010111110010101110011010001001100000110000101111100101011100110100010010000011100001011111001010111001101000100000000111000010111110010101110011010001000000001110000101111100101011100110100010000000001011111001010111001101000100111100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b100010100001100000100000011111110101000001000101000011000001000000111111101000000110001010000110000010000001111111010000011100010100001100000100000011111110000001111000101000011000001000000111111100000011110001010000110000010000001111110000000010100001100000100000011111110101000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b010011001110111010010110001101111011000000100110011101110100101100011011110100000101001100111011101001011000110111100000001010011001110111010010110001101111000001010100110011101110100101100011011100000010101001100111011101001011000110110000010011001110111010010110001101111011000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b010110110010010001110000101111100101000000101101100100100011100001011111001000000101011011001001000111000010111110010000011010110110010010001110000101111100000000110101101100100100011100001011111000000101101011011001001000111000010111110000010110110010010001110000101111100101000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b011100110100010011110001010000110000000000111001101000100111100010100001100000000101110011010001001111000101000011000000001011100110100010011110001010000110000001010111001101000100111100010100001100000010101110011010001001111000101000010000011100110100010011110001010000110000000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b010000001111111010101001100111011101000000100000011111110101010011001110111000000001000000111111101010100110011101110000000010000001111111010101001100111011000000000100000011111110101010011001110100000000001000000111111101010100110011100000010000001111111010101001100111011101000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b001011000110111101101011011001001000000000010110001101111011010110110010010000000100101100011011110110101101100100100000001001011000110111101101011011001001000001010010110001101111011010110110010000000110100101100011011110110101101100100000001011000110111101101011011001001000100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b111000010111110010101110011010001001000001110000101111100101011100110100010000000011100001011111001010111001101000100000000111000010111110010101110011010001000000001110000101111100101011100110100000000100011100001011111001010111001101000000011000010111110010101110011010001001100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b111000101000011000001000000111111101000001110001010000110000010000001111111000000111100010100001100000100000011111110000001111000101000011000001000000111111000000011110001010000110000010000001111100000100111100010100001100000100000011110000011000101000011000001000000111111101000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b010100110011101110100101100011011110000000101001100111011101001011000110111100000101010011001110111010010110001101110000001010100110011101110100101100011011000001010101001100111011101001011000110100000110101010011001110111010010110001100000010100110011101110100101100011011110100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b110101101100100100011100001011111001000001101011011001001000111000010111110000000011010110110010010001110000101111100000010110101101100100100011100001011111000001101101011011001001000111000010111100000111011010110110010010001110000101110000010101101100100100011100001011111001000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b010111001101000100111100010100001100000000101110011010001001111000101000011000000101011100110100010011110001010000110000001010111001101000100111100010100001000000010101110011010001001111000101000000000100101011100110100010011110001010000000010111001101000100111100010100001100000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b000100000011111110101010011001110111000000001000000111111101010100110011101100000000010000001111111010101001100111010000000000100000011111110101010011001110000001000001000000111111101010100110011100000110000010000001111111010101001100110000000100000011111110101010011001110111000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b010010110001101111011010110110010010000000100101100011011110110101101100100100000101001011000110111101101011011001000000011010010110001101111011010110110010000001110100101100011011110110101101100100000011101001011000110111101101011011000000010010110001101111011010110110010010000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b001110000101111100101011100110100010000000011100001011111001010111001101000100000000111000010111110010101110011010000000010001110000101111100101011100110100000000100011100001011111001010111001101000000001000111000010111110010101110011010000001110000101111100101011100110100010000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b011110001010000110000010000001111111000000111100010100001100000100000011111100000001111000101000011000001000000111110000010011110001010000110000010000001111000000100111100010100001100000100000011100000001001111000101000011000001000000110000011110001010000110000010000001111111000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b010101001100111011101001011000110111000000101010011001110111010010110001101100000101010100110011101110100101100011010000011010101001100111011101001011000110000001110101010011001110111010010110001100000111101010100110011101110100101100010000010101001100111011101001011000110111100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b101101011011001001000111000010111110000001011010110110010010001110000101111100000110110101101100100100011100001011110000011101101011011001001000111000010111000001111011010110110010010001110000101100000011110110101101100100100011100001010000001101011011001001000111000010111110000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b010101110011010001001111000101000011000000101011100110100010011110001010000100000001010111001101000100111100010100000000010010101110011010001001111000101000000001100101011100110100010011110001010000000111001010111001101000100111100010100000010101110011010001001111000101000011000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b000001000000111111101010100110011101000000000010000001111111010101001100111000000100000100000011111110101010011001110000011000001000000111111101010100110011000000110000010000001111111010101001100100000001100000100000011111110101010011000000000001000000111111101010100110011101100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b110100101100011011110110101101100100000001101001011000110111101101011011001000000111010010110001101111011010110110010000001110100101100011011110110101101100000001011101001011000110111101101011011000000110111010010110001101111011010110110000010100101100011011110110101101100100100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b100011100001011111001010111001101000000001000111000010111110010101110011010000000010001110000101111100101011100110100000000100011100001011111001010111001101000001001000111000010111110010101110011000000010010001110000101111100101011100110000000011100001011111001010111001101000100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b100111100010100001100000100000011111000001001111000101000011000001000000111100000010011110001010000110000010000001110000000100111100010100001100000100000011000000001001111000101000011000001000000100000100010011110001010000110000010000000000000111100010100001100000100000011111100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b110101010011001110111010010110001101000001101010100110011101110100101100011000000111010101001100111011101001011000110000011110101010011001110111010010110001000001111101010100110011101110100101100000000111111010101001100111011101001011000000010101010011001110111010010110001101100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b111011010110110010010001110000101111000001110110101101100100100011100001011100000111101101011011001001000111000010110000001111011010110110010010001110000101000001011110110101101100100100011100001000000110111101101011011001001000111000010000011011010110110010010001110000101111100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b100101011100110100010011110001010000000001001010111001101000100111100010100000000110010101110011010001001111000101000000011100101011100110100010011110001010000001111001010111001101000100111100010100000111110010101110011010001001111000100000000101011100110100010011110001010000100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b110000010000001111111010101001100111000001100000100000011111110101010011001100000011000001000000111111101010100110010000000110000010000001111111010101001100000000001100000100000011111110101010011000000000011000001000000111111101010100110000010000010000001111111010101001100111000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b011101001011000110111101101011011001000000111010010110001101111011010110110000000101110100101100011011110110101101100000011011101001011000110111101101011011000001110111010010110001101111011010110100000011101110100101100011011110110101100000011101001011000110111101101011011001000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b001000111000010111110010101110011010000000010001110000101111100101011100110100000100100011100001011111001010111001100000001001000111000010111110010101110011000000010010001110000101111100101011100100000100100100011100001011111001010111000000001000111000010111110010101110011010000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b001001111000101000011000001000000111000000010011110001010000110000010000001100000000100111100010100001100000100000010000010001001111000101000011000001000000000000100010011110001010000110000010000000000101000100111100010100001100000100000000001001111000101000011000001000000111100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b111101010100110011101110100101100011000001111010101001100111011101001011000100000111110101010011001110111010010110000000011111101010100110011101110100101100000001111111010101001100111011101001011000000011111110101010011001110111010010110000011101010100110011101110100101100011000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b011110110101101100100100011100001011000000111101101011011001001000111000010100000101111011010110110010010001110000100000011011110110101101100100100011100001000000110111101101011011001001000111000000000001101111011010110110010010001110000000011110110101101100100100011100001011100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b111001010111001101000100111100010100000001110010101110011010001001111000101000000111100101011100110100010011110001010000011111001010111001101000100111100010000000111110010101110011010001001111000100000101111100101011100110100010011110000000011001010111001101000100111100010100000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b001100000100000011111110101010011001000000011000001000000111111101010100110000000000110000010000001111111010101001100000000001100000100000011111110101010011000001000011000001000000111111101010100100000010000110000010000001111111010101000000001100000100000011111110101010011001100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b110111010010110001101111011010110110000001101110100101100011011110110101101100000111011101001011000110111101101011010000001110111010010110001101111011010110000000011101110100101100011011110110101100000100111011101001011000110111101101010000010111010010110001101111011010110110000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b010010001110000101111100101011100110000000100100011100001011111001010111001100000001001000111000010111110010101110010000010010010001110000101111100101011100000001100100100011100001011111001010111000000011001001000111000010111110010101110000010010001110000101111100101011100110100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b100010011110001010000110000010000001000001000100111100010100001100000100000000000010001001111000101000011000001000000000010100010011110001010000110000010000000001101000100111100010100001100000100000000011010001001111000101000011000001000000000010011110001010000110000010000001100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b111111010101001100111011101001011000000001111110101010011001110111010010110000000111111101010100110011101110100101100000001111111010101001100111011101001011000000011111110101010011001110111010010100000000111111101010100110011101110100100000011111010101001100111011101001011000100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b110111101101011011001001000111000010000001101111011010110110010010001110000100000011011110110101101100100100011100000000000110111101101011011001001000111000000000001101111011010110110010010001110000000100011011110110101101100100100011100000010111101101011011001001000111000010100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b111110010101110011010001001111000101000001111100101011100110100010011110001000000011111001010111001101000100111100010000010111110010101110011010001001111000000000101111100101011100110100010011110000000001011111001010111001101000100111100000011110010101110011010001001111000101000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b000011000001000000111111101010100110000000000110000010000001111111010101001100000100001100000100000011111110101010010000001000011000001000000111111101010100000001010000110000010000001111111010101000000010100001100000100000011111110101010000000011000001000000111111101010100110000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b011101110100101100011011110110101101000000111011101001011000110111101101011000000001110111010010110001101111011010110000010011101110100101100011011110110101000001100111011101001011000110111101101000000011001110111010010110001101111011010000011101110100101100011011110110101101100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b100100100011100001011111001010111001000001001001000111000010111110010101110000000110010010001110000101111100101011100000001100100100011100001011111001010111000001011001001000111000010111110010101100000110110010010001110000101111100101010000000100100011100001011111001010111001100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b101000100111100010100001100000100000000001010001001111000101000011000001000000000110100010011110001010000110000010000000001101000100111100010100001100000100000000011010001001111000101000011000001000000100110100010011110001010000110000010000001000100111100010100001100000100000000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b011111110101010011001110111010010110000000111111101010100110011101110100101100000001111111010101001100111011101001010000000011111110101010011001110111010010000000000111111101010100110011101110100100000000001111111010101001100111011101000000011111110101010011001110111010010110000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b001101111011010110110010010001110000000000011011110110101101100100100011100000000000110111101101011011001001000111000000010001101111011010110110010010001110000001100011011110110101101100100100011100000011000110111101101011011001001000110000001101111011010110110010010001110000100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b101111100101011100110100010011110001000001011111001010111001101000100111100000000010111110010101110011010001001111000000000101111100101011100110100010011110000000001011111001010111001101000100111100000000010111110010101110011010001001110000001111100101011100110100010011110001000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b010000110000010000001111111010101001000000100001100000100000011111110101010000000101000011000001000000111111101010100000001010000110000010000001111111010101000000010100001100000100000011111110101000000000101000011000001000000111111101010000010000110000010000001111111010101001100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b100111011101001011000110111101101011000001001110111010010110001101111011010100000110011101110100101100011011110110100000001100111011101001011000110111101101000000011001110111010010110001101111011000000100110011101110100101100011011110110000000111011101001011000110111101101011000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b011001001000111000010111110010101110000000110010010001110000101111100101011100000101100100100011100001011111001010110000011011001001000111000010111110010101000000110110010010001110000101111100101000000101101100100100011100001011111001010000011001001000111000010111110010101110000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b011010001001111000101000011000001000000000110100010011110001010000110000010000000001101000100111100010100001100000100000010011010001001111000101000011000001000001100110100010011110001010000110000000000111001101000100111100010100001100000000011010001001111000101000011000001000000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b000111111101010100110011101110100101000000001111111010101001100111011101001000000000011111110101010011001110111010010000000000111111101010100110011101110100000000000001111111010101001100111011101000000100000011111110101010011001110111010000000111111101010100110011101110100101100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b100011011110110101101100100100011100000001000110111101101011011001001000111000000110001101111011010110110010010001110000001100011011110110101101100100100011000001011000110111101101011011001001000100000010110001101111011010110110010010000000000011011110110101101100100100011100000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b001011111001010111001101000100111100000000010111110010101110011010001001111000000000101111100101011100110100010011110000000001011111001010111001101000100111000001000010111110010101110011010001001100000110000101111100101011100110100010010000001011111001010111001101000100111100000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b010100001100000100000011111110101010000000101000011000001000000111111101010100000001010000110000010000001111111010100000000010100001100000100000011111110101000001000101000011000001000000111111101000000110001010000110000010000001111111010000010100001100000100000011111110101010000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b011001110111010010110001101111011010000000110011101110100101100011011110110100000001100111011101001011000110111101100000010011001110111010010110001101111011000000100110011101110100101100011011110100000101001100111011101001011000110111100000011001110111010010110001101111011010100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b110110010010001110000101111100101011000001101100100100011100001011111001010100000011011001001000111000010111110010100000010110110010010001110000101111100101000000101101100100100011100001011111001000000101011011001001000111000010111110010000010110010010001110000101111100101011100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b100110100010011110001010000110000010000001001101000100111100010100001100000100000110011010001001111000101000011000000000011100110100010011110001010000110000000000111001101000100111100010100001100000000101110011010001001111000101000011000000000110100010011110001010000110000010000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b000001111111010101001100111011101001000000000011111110101010011001110111010000000000000111111101010100110011101110100000010000001111111010101001100111011101000000100000011111110101010011001110111000000001000000111111101010100110011101110000000001111111010101001100111011101001000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b011000110111101101011011001001000111000000110001101111011010110110010010001100000101100011011110110101101100100100010000001011000110111101101011011001001000000000010110001101111011010110110010010000000100101100011011110110101101100100100000011000110111101101011011001001000111000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b000010111110010101110011010001001111000000000101111100101011100110100010011100000100001011111001010111001101000100110000011000010111110010101110011010001001000001110000101111100101011100110100010000000011100001011111001010111001101000100000000010111110010101110011010001001111000000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b000101000011000001000000111111101010000000001010000110000010000001111111010100000100010100001100000100000011111110100000011000101000011000001000000111111101000001110001010000110000010000001111111000000111100010100001100000100000011111110000000101000011000001000000111111101010100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b100110011101110100101100011011110110000001001100111011101001011000110111101100000010011001110111010010110001101111010000010100110011101110100101100011011110000000101001100111011101001011000110111100000101010011001110111010010110001101110000000110011101110100101100011011110110100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b101101100100100011100001011111001010000001011011001001000111000010111110010100000010110110010010001110000101111100100000010101101100100100011100001011111001000001101011011001001000111000010111110000000011010110110010010001110000101111100000001101100100100011100001011111001010100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);

#5 CK=0;
#5 LFSR=247'b111001101000100111100010100001100000000001110011010001001111000101000011000000000011100110100010011110001010000110000000010111001101000100111100010100001100000000101110011010001001111000101000011000000101011100110100010011110001010000110000011001101000100111100010100001100000100000;
#5 CK=1;
$fwrite(f, "%b\n", TEST_OUT);


      $fclose(f);
   end


endmodule // nm_testbench
